// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, the Altera Quartus Prime License Agreement,
// the Altera MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Altera and sold by Altera or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// Generated by Quartus Prime Version 15.1.1 Build 189 12/02/2015 SJ Lite Edition
// Created on Mon Nov 14 05:32:26 2016

// synthesis message_off 10175

`timescale 1ns/1ns

module nothing2 (
    reset,clock,x,
    z,t,fstate);

    input reset;
    input clock;
    input x;
    tri0 reset;
    tri0 x;
    output z;
    output t;
    reg z;
    reg t;
    output reg [2:0] fstate;
    reg [2:0] reg_fstate;
    parameter xxx=0,qqq=1,state1=2;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or x)
    begin
        if (reset) begin
            reg_fstate <= xxx;
            z <= 1'b0;
            t <= 1'b0;
        end
        else begin
            z <= 1'b0;
            t <= 1'b0;
            case (fstate)
                xxx: begin
                    reg_fstate <= qqq;

                    if (x)
                        t <= 1'b1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        t <= 1'b0;
                end
                qqq: begin
                    if (x)
                        reg_fstate <= state1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= qqq;

                    z <= 1'b1;
                end
                state1: begin
                    if (x)
                        reg_fstate <= xxx;
                    else
                        reg_fstate <= state1;
                end
                default: begin
                    z <= 1'bx;
                    t <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // nothing2
