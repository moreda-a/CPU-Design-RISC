reg8_SP_inst : reg8_SP PORT MAP (
		aclr	 => aclr_sig,
		clock	 => clock_sig,
		cnt_en	 => cnt_en_sig,
		sset	 => sset_sig,
		updown	 => updown_sig,
		q	 => q_sig
	);
