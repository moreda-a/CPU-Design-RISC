-- Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, the Altera Quartus Prime License Agreement,
-- the Altera MegaCore Function License Agreement, or other 
-- applicable license agreement, including, without limitation, 
-- that your use is for the sole purpose of programming logic 
-- devices manufactured by Altera and sold by Altera or its 
-- authorized distributors.  Please refer to the applicable 
-- agreement for further details.

-- Generated by Quartus Prime Version 15.1.1 Build 189 12/02/2015 SJ Lite Edition
-- Created on Mon Nov 14 05:03:14 2016

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY nothing2 IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        x : IN STD_LOGIC := '0';
        z : OUT STD_LOGIC;
        t : OUT STD_LOGIC
    );
END nothing2;

ARCHITECTURE BEHAVIOR OF nothing2 IS
    TYPE type_fstate IS (qqq,state3,xxx);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,x)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= xxx;
            z <= '0';
            t <= '0';
        ELSE
            z <= '0';
            t <= '0';
            CASE fstate IS
                WHEN qqq =>
                    reg_fstate <= state3;

                    z <= '1';
                WHEN state3 =>
                    reg_fstate <= xxx;
                WHEN xxx =>
                    reg_fstate <= qqq;

                    IF ((x = '1')) THEN
                        t <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        t <= '0';
                    END IF;
                WHEN OTHERS => 
                    z <= 'X';
                    t <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
